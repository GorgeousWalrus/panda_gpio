
`define GPIO_DIR 0
`define GPIO_VAL 1
`define GPIO_INV 2
`define GPIO_INT_EN 3
`define GPIO_INT_T 4

`define GPIO_INT_T_RISE 1'b0
`define GPIO_INT_T_EDGE 1'b1